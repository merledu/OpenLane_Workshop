VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO manual_macro_placement_test
  CLASS BLOCK ;
  FOREIGN manual_macro_placement_test ;
  ORIGIN 0.000 0.000 ;
  SIZE 312.060 BY 322.780 ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 61.240 312.060 61.840 ;
    END
  END clk2
  PIN p1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 318.780 34.870 322.780 ;
    END
  END p1
  PIN p2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 167.320 312.060 167.920 ;
    END
  END p2
  PIN rst1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END rst1
  PIN rst2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 275.440 312.060 276.040 ;
    END
  END rst2
  PIN x1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END x1[0]
  PIN x1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 318.780 294.310 322.780 ;
    END
  END x1[10]
  PIN x1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END x1[11]
  PIN x1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END x1[12]
  PIN x1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 318.780 21.070 322.780 ;
    END
  END x1[13]
  PIN x1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END x1[14]
  PIN x1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 104.080 312.060 104.680 ;
    END
  END x1[15]
  PIN x1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 318.780 63.850 322.780 ;
    END
  END x1[16]
  PIN x1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END x1[17]
  PIN x1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 318.780 265.330 322.780 ;
    END
  END x1[18]
  PIN x1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END x1[19]
  PIN x1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END x1[1]
  PIN x1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 318.780 207.370 322.780 ;
    END
  END x1[20]
  PIN x1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END x1[21]
  PIN x1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END x1[22]
  PIN x1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 318.780 5.890 322.780 ;
    END
  END x1[23]
  PIN x1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END x1[24]
  PIN x1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END x1[25]
  PIN x1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END x1[26]
  PIN x1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 318.780 280.510 322.780 ;
    END
  END x1[27]
  PIN x1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 318.780 308.110 322.780 ;
    END
  END x1[28]
  PIN x1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 83.680 312.060 84.280 ;
    END
  END x1[29]
  PIN x1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 253.000 312.060 253.600 ;
    END
  END x1[2]
  PIN x1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 318.780 178.390 322.780 ;
    END
  END x1[30]
  PIN x1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END x1[31]
  PIN x1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 126.520 312.060 127.120 ;
    END
  END x1[3]
  PIN x1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END x1[4]
  PIN x1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 318.780 164.590 322.780 ;
    END
  END x1[5]
  PIN x1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END x1[6]
  PIN x1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 318.780 236.350 322.780 ;
    END
  END x1[7]
  PIN x1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END x1[8]
  PIN x1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 40.840 312.060 41.440 ;
    END
  END x1[9]
  PIN x2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END x2[0]
  PIN x2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 318.780 121.810 322.780 ;
    END
  END x2[10]
  PIN x2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END x2[11]
  PIN x2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END x2[12]
  PIN x2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 18.400 312.060 19.000 ;
    END
  END x2[13]
  PIN x2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 318.780 193.570 322.780 ;
    END
  END x2[14]
  PIN x2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 318.780 150.790 322.780 ;
    END
  END x2[15]
  PIN x2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 318.780 92.830 322.780 ;
    END
  END x2[16]
  PIN x2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END x2[17]
  PIN x2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 318.780 106.630 322.780 ;
    END
  END x2[18]
  PIN x2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 295.840 312.060 296.440 ;
    END
  END x2[19]
  PIN x2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END x2[1]
  PIN x2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END x2[20]
  PIN x2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END x2[21]
  PIN x2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 210.160 312.060 210.760 ;
    END
  END x2[22]
  PIN x2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END x2[23]
  PIN x2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 318.780 251.530 322.780 ;
    END
  END x2[24]
  PIN x2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 318.780 222.550 322.780 ;
    END
  END x2[25]
  PIN x2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 189.760 312.060 190.360 ;
    END
  END x2[26]
  PIN x2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END x2[27]
  PIN x2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END x2[28]
  PIN x2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END x2[29]
  PIN x2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 318.780 77.650 322.780 ;
    END
  END x2[2]
  PIN x2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END x2[30]
  PIN x2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 146.920 312.060 147.520 ;
    END
  END x2[31]
  PIN x2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END x2[3]
  PIN x2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.060 232.600 312.060 233.200 ;
    END
  END x2[4]
  PIN x2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END x2[5]
  PIN x2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END x2[6]
  PIN x2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 318.780 135.610 322.780 ;
    END
  END x2[7]
  PIN x2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END x2[8]
  PIN x2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END x2[9]
  PIN y1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 318.780 48.670 322.780 ;
    END
  END y1
  PIN y2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END y2
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 154.720 10.640 156.320 310.320 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 274.720 10.640 276.320 158.470 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 244.720 10.640 246.320 158.470 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 214.720 10.640 216.320 158.470 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.720 10.640 186.320 158.470 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 124.720 10.640 126.320 158.470 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 94.720 10.640 96.320 158.470 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 64.720 10.640 66.320 158.470 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 34.720 10.640 36.320 158.470 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 306.360 181.270 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 306.360 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 139.720 10.640 141.320 310.320 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 289.720 10.640 291.320 158.470 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 259.720 10.640 261.320 158.470 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 229.720 10.640 231.320 158.470 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 199.720 10.640 201.320 158.470 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 169.720 10.640 171.320 158.470 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 109.720 10.640 111.320 158.470 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 79.720 10.640 81.320 158.470 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.720 10.640 51.320 158.470 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 19.720 10.640 21.320 158.470 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 306.360 257.860 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 306.360 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 7.045 11.305 304.835 311.015 ;
      LAYER met1 ;
        RECT 2.830 9.560 308.130 312.420 ;
      LAYER met2 ;
        RECT 2.860 318.500 5.330 318.780 ;
        RECT 6.170 318.500 20.510 318.780 ;
        RECT 21.350 318.500 34.310 318.780 ;
        RECT 35.150 318.500 48.110 318.780 ;
        RECT 48.950 318.500 63.290 318.780 ;
        RECT 64.130 318.500 77.090 318.780 ;
        RECT 77.930 318.500 92.270 318.780 ;
        RECT 93.110 318.500 106.070 318.780 ;
        RECT 106.910 318.500 121.250 318.780 ;
        RECT 122.090 318.500 135.050 318.780 ;
        RECT 135.890 318.500 150.230 318.780 ;
        RECT 151.070 318.500 164.030 318.780 ;
        RECT 164.870 318.500 177.830 318.780 ;
        RECT 178.670 318.500 193.010 318.780 ;
        RECT 193.850 318.500 206.810 318.780 ;
        RECT 207.650 318.500 221.990 318.780 ;
        RECT 222.830 318.500 235.790 318.780 ;
        RECT 236.630 318.500 250.970 318.780 ;
        RECT 251.810 318.500 264.770 318.780 ;
        RECT 265.610 318.500 279.950 318.780 ;
        RECT 280.790 318.500 293.750 318.780 ;
        RECT 294.590 318.500 307.550 318.780 ;
        RECT 2.860 4.280 308.100 318.500 ;
        RECT 3.410 4.000 16.370 4.280 ;
        RECT 17.210 4.000 30.170 4.280 ;
        RECT 31.010 4.000 45.350 4.280 ;
        RECT 46.190 4.000 59.150 4.280 ;
        RECT 59.990 4.000 74.330 4.280 ;
        RECT 75.170 4.000 88.130 4.280 ;
        RECT 88.970 4.000 103.310 4.280 ;
        RECT 104.150 4.000 117.110 4.280 ;
        RECT 117.950 4.000 132.290 4.280 ;
        RECT 133.130 4.000 146.090 4.280 ;
        RECT 146.930 4.000 159.890 4.280 ;
        RECT 160.730 4.000 175.070 4.280 ;
        RECT 175.910 4.000 188.870 4.280 ;
        RECT 189.710 4.000 204.050 4.280 ;
        RECT 204.890 4.000 217.850 4.280 ;
        RECT 218.690 4.000 233.030 4.280 ;
        RECT 233.870 4.000 246.830 4.280 ;
        RECT 247.670 4.000 262.010 4.280 ;
        RECT 262.850 4.000 275.810 4.280 ;
        RECT 276.650 4.000 289.610 4.280 ;
        RECT 290.450 4.000 304.790 4.280 ;
        RECT 305.630 4.000 308.100 4.280 ;
      LAYER met3 ;
        RECT 4.000 302.960 308.060 311.945 ;
        RECT 4.400 301.560 308.060 302.960 ;
        RECT 4.000 296.840 308.060 301.560 ;
        RECT 4.000 295.440 307.660 296.840 ;
        RECT 4.000 280.520 308.060 295.440 ;
        RECT 4.400 279.120 308.060 280.520 ;
        RECT 4.000 276.440 308.060 279.120 ;
        RECT 4.000 275.040 307.660 276.440 ;
        RECT 4.000 260.120 308.060 275.040 ;
        RECT 4.400 258.720 308.060 260.120 ;
        RECT 4.000 254.000 308.060 258.720 ;
        RECT 4.000 252.600 307.660 254.000 ;
        RECT 4.000 237.680 308.060 252.600 ;
        RECT 4.400 236.280 308.060 237.680 ;
        RECT 4.000 233.600 308.060 236.280 ;
        RECT 4.000 232.200 307.660 233.600 ;
        RECT 4.000 217.280 308.060 232.200 ;
        RECT 4.400 215.880 308.060 217.280 ;
        RECT 4.000 211.160 308.060 215.880 ;
        RECT 4.000 209.760 307.660 211.160 ;
        RECT 4.000 194.840 308.060 209.760 ;
        RECT 4.400 193.440 308.060 194.840 ;
        RECT 4.000 190.760 308.060 193.440 ;
        RECT 4.000 189.360 307.660 190.760 ;
        RECT 4.000 174.440 308.060 189.360 ;
        RECT 4.400 173.040 308.060 174.440 ;
        RECT 4.000 168.320 308.060 173.040 ;
        RECT 4.000 166.920 307.660 168.320 ;
        RECT 4.000 154.040 308.060 166.920 ;
        RECT 4.400 152.640 308.060 154.040 ;
        RECT 4.000 147.920 308.060 152.640 ;
        RECT 4.000 146.520 307.660 147.920 ;
        RECT 4.000 131.600 308.060 146.520 ;
        RECT 4.400 130.200 308.060 131.600 ;
        RECT 4.000 127.520 308.060 130.200 ;
        RECT 4.000 126.120 307.660 127.520 ;
        RECT 4.000 111.200 308.060 126.120 ;
        RECT 4.400 109.800 308.060 111.200 ;
        RECT 4.000 105.080 308.060 109.800 ;
        RECT 4.000 103.680 307.660 105.080 ;
        RECT 4.000 88.760 308.060 103.680 ;
        RECT 4.400 87.360 308.060 88.760 ;
        RECT 4.000 84.680 308.060 87.360 ;
        RECT 4.000 83.280 307.660 84.680 ;
        RECT 4.000 68.360 308.060 83.280 ;
        RECT 4.400 66.960 308.060 68.360 ;
        RECT 4.000 62.240 308.060 66.960 ;
        RECT 4.000 60.840 307.660 62.240 ;
        RECT 4.000 45.920 308.060 60.840 ;
        RECT 4.400 44.520 308.060 45.920 ;
        RECT 4.000 41.840 308.060 44.520 ;
        RECT 4.000 40.440 307.660 41.840 ;
        RECT 4.000 25.520 308.060 40.440 ;
        RECT 4.400 24.120 308.060 25.520 ;
        RECT 4.000 19.400 308.060 24.120 ;
        RECT 4.000 18.000 307.660 19.400 ;
        RECT 4.000 9.015 308.060 18.000 ;
      LAYER met4 ;
        RECT 6.735 310.720 299.130 311.945 ;
        RECT 6.735 158.870 139.320 310.720 ;
        RECT 6.735 10.240 19.320 158.870 ;
        RECT 21.720 10.240 34.320 158.870 ;
        RECT 36.720 10.240 49.320 158.870 ;
        RECT 51.720 10.240 64.320 158.870 ;
        RECT 66.720 10.240 79.320 158.870 ;
        RECT 81.720 10.240 94.320 158.870 ;
        RECT 96.720 10.240 109.320 158.870 ;
        RECT 111.720 10.240 124.320 158.870 ;
        RECT 126.720 10.240 139.320 158.870 ;
        RECT 141.720 10.240 154.320 310.720 ;
        RECT 156.720 158.870 299.130 310.720 ;
        RECT 156.720 10.240 169.320 158.870 ;
        RECT 171.720 10.240 184.320 158.870 ;
        RECT 186.720 10.240 199.320 158.870 ;
        RECT 201.720 10.240 214.320 158.870 ;
        RECT 216.720 10.240 229.320 158.870 ;
        RECT 231.720 10.240 244.320 158.870 ;
        RECT 246.720 10.240 259.320 158.870 ;
        RECT 261.720 10.240 274.320 158.870 ;
        RECT 276.720 10.240 289.320 158.870 ;
        RECT 291.720 10.240 299.130 158.870 ;
        RECT 6.735 9.015 299.130 10.240 ;
      LAYER met5 ;
        RECT 7.940 259.460 299.340 274.500 ;
        RECT 7.940 215.100 299.340 254.660 ;
  END
END manual_macro_placement_test
END LIBRARY

